module IF_Stage (input clk, rst, output[31:0] PC, Instruction);

endmodule