module tb();
    MIPS(.clk(clk), .rst(rst));

    wire clk = 0, rst = 1;
    

endmodule