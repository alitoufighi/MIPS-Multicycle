`timescale 1ns/1ns
module tb();
  reg clk                     = 1, rst = 1;
  wire [17:0]s;
  assign s                    = {14'b0, rst, 3'b0};
  
  wire [15:0] SRAM_DQ;
  wire [17:0] SRAM_ADDR;
  wire SRAM_WE_N;

	MIPS mips(
			.CLOCK_50(clk),
			.SW(s), 
		   	.SRAM_DQ(SRAM_DQ),           // SRAM Data bus
		    .SRAM_ADDR(SRAM_ADDR),    // SRAM Addr bus
			.SRAM_WE_N(SRAM_WE_N)          // SRAM write enable
	);

	SRAM sram(clk, rst, SRAM_DQ, SRAM_ADDR, SRAM_WE_N);

	initial begin
		#20 rst               =~rst;

		repeat(900)#10 clk    =~clk;
	end
    
endmodule

