module MEM_Stage_reg(input clk, rst, input[31:0] PC_in, output reg[31:0] PC);

endmodule